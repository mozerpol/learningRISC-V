`define EQ 3'b000
`define NE 3'b001
`define LT 3'b010
`define GE 3'b011 
`define LTU 3'b100
`define GEU 3'b101