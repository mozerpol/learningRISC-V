library ieee;
   use ieee.std_logic_1164.all;
   use ieee.numeric_std.all;
   use ieee.std_logic_unsigned.all;
library std;
  use std.env.all;

entity main_tb is
end main_tb;

architecture tb of main_tb is

   component main is
   port (
      i_rst                : in std_logic;
      i_clk                : in std_logic;
      i_instruction_read   : in std_logic_vector(31 downto 0);
      o_instruction_write  : out std_logic_vector(31 downto 0);
      o_addr_read          : out std_logic_vector(7 downto 0);
      o_addr_write         : out std_logic_vector(7 downto 0);
      o_write_enable       : out std_logic
   );
   end component main;

   signal rst_tb              : std_logic;
   signal clk_tb              : std_logic;
   signal instruction_read_tb      : std_logic_vector(31 downto 0);
   signal instruction_write_tb    : std_logic_vector(31 downto 0);
   signal addr_read_tb    : std_logic_vector(7 downto 0);
   signal addr_write_tb   : std_logic_vector(7 downto 0);
   signal write_enable_tb : std_logic;

begin

   inst_main : component main
   port map (
      i_rst                => rst_tb,
      i_clk                => clk_tb,
      i_instruction_read        => instruction_read_tb,
      o_instruction_write      => instruction_write_tb,
      o_addr_read          => addr_read_tb,
      o_addr_write         => addr_write_tb,
      o_write_enable       => write_enable_tb
   );




end architecture tb;
