library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
   use ieee.numeric_std.all;
library rysy_pkg;
   use rysy_pkg.rysyPkg.all;
library imm_mux_lib;
   use imm_mux_lib.all;
   use imm_mux_lib.imm_mux_pkg.all;

entity imm_mux is
   port (
   );
end entity imm_mux;

architecture rtl of imm_mux is

begin

   p_imm_mux : process(all)
   begin
   end process p_imm_mux;

end architecture rtl;
