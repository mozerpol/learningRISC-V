library ieee;
   use ieee.std_logic_1164.all;
   use ieee.numeric_std.all;
   use ieee.std_logic_unsigned.all;
   
package rysy_pkg is
   -- constant C_NAME : std_logic_vector(N downto M) := "X";
end;
 
package body rysy_pkg is
 
end package body;
