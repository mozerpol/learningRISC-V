`define	INST_OLD 2'b00
`define INST_NOP 2'b01
`define INST_MEM 2'b10