library ieee;
   use ieee.std_logic_1164.all;
   use IEEE.std_logic_unsigned.all;
   use IEEE.math_real.all;

 package alu_mux_1_pkg is
    -- constant C_NAME : std_logic_vector(N downto M) := "X";
    constant C_RS1_DATA : std_logic := '0';
    constant C_PC_ADDR  : std_logic := '1';

 end;

 package body alu_mux_1_pkg is

 end package body;
