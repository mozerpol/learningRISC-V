library ieee;
   use ieee.std_logic_1164.all;
   use ieee.numeric_std.all;
   use ieee.std_logic_unsigned.all;
library rysy_pkg;
   use rysy_pkg.rysyPkg.all;

entity alu1_mux_tb is
end alu1_mux_tb;

architecture tb of alu1_mux_tb is
begin

end architecture tb;
