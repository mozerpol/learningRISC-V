--------------------------------------------------------------------------------
-- File          : riscpol_pkg.vhdl
-- Author        : mozerpol
--------------------------------------------------------------------------------
-- Description   : Package with RAM and ROM size settings and addresses, which
-- control access to external peripherals, e.g. at what address is access to
-- GPIO or TIMER.
--------------------------------------------------------------------------------
-- License       : MIT 2022 mozerpol
--------------------------------------------------------------------------------


library ieee;
   use ieee.std_logic_1164.all;


package riscpol_pkg is


   constant C_CLK_PERIOD      : time    := 20 ns; -- Constant needed only for  50000000
   constant C_FREQUENCY_MHZ   : positive := positive(1.0/(real(C_CLK_PERIOD/ns)/1000000000.0));
   -- test purposes.
   constant C_RAM_BYTE_WIDTH  : natural := 8;    -- For RAM purposes, don't
   -- touch, constant is generated by Quartus, as a part of template
   -- "Byte-enabled Simple Dual Port RAM".
   constant C_RAM_BYTES       : natural := 4;    -- As above
   constant C_RAM_LENGTH      : integer := 64;   -- RAM size in
   -- peripherals/ram.vhdl file. If you want to have more memory for data (for 
   -- instructions is C_ROM_LENGTH) change this value.
   constant C_ROM_LENGTH      : integer := 1024; -- Instruction memory size that
   -- changes the size of C_CODE array in instruction_memory_design.vhdl file.
   -- Must be greater than or equal to the number of instructions and a power of
   -- number 2.
   constant C_MMIO_ADDR_GPIO  : integer := 64;   -- At what address is access to
   -- GPIO. To know more about MMIO take a look at Wikipedia.
   constant C_MMIO_ADDR_CNT_8_BIT : integer := 63;   --
   constant C_MMIO_ADDR_UART : integer := 62;   --
   --constant C_MMIO_ADDR_UART_DATA : integer := 61;   --
   
   constant C_COUNTER_8BIT_VALUE : integer := 512;   -- Up to what value should 
   -- the counter 8 bit count?
   
   constant C_NUMBER_OF_GPIO : integer := 8;   -- 
   
   constant C_BAUD : positive := 115200;   -- 

   -- Type for General-Purpose Register
   type t_gpr  is array(0 to 31) of std_logic_vector(31 downto 0);
   --  Build up 2D array to hold the data memory (ram.vhd)
   type word_t is array (0 to C_RAM_BYTES-1) of std_logic_vector(C_RAM_BYTE_WIDTH-1 downto 0);
   type ram_t is array (0 to C_RAM_LENGTH - 1) of word_t;


end;


package body riscpol_pkg is


end package body;
