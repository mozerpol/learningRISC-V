library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
   use ieee.numeric_std.all;
library rysy_pkg;
   use rysy_pkg.rysyPkg.all;
library mem_addr_sel_lib;
   use mem_addr_sel_lib.all;
   use mem_addr_sel_lib.mem_addr_sel_pkg.all;

entity mem_addr_sel is
   port (
   );
end entity mem_addr_sel;

architecture rtl of mem_addr_sel is

begin

   p_mem_addr_sel : process(all)
   begin
   end process p_mem_addr_sel;

end architecture rtl;
