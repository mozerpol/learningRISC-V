library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
   use ieee.numeric_std.all;
library rysy_pkg;
   use rysy_pkg.rysyPkg.all;


entity select_rd_design is
   );
end entity select_rd_design;

architecture rtl of select_rd_design is

begin

end architecture rtl;
