`timescale 100ns / 10ns

// SB, SH, ... are S-type instructions, storage instructions.

`define SB  3'b000
`define SH  3'b001
`define SW  3'b010
`define SBU 3'b011
`define SHU 3'b100

module sel_type(
  input [2:0] sel_type_input,
  output [2:0] sel_type_output
);

	assign sel_type_output = sel_type_input;

endmodule
