library ieee;
   use ieee.std_logic_1164.all;
   use IEEE.std_logic_unsigned.all;
   use IEEE.math_real.all;

 package mmio_pkg is

 end;

 package body mmio_pkg is

 end package body;
