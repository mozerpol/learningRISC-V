library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
   use ieee.numeric_std.all;
library memory_management_lib;
   use memory_management_lib.all;
   use memory_management_lib.memory_management_pkg.all;

entity memory_management is
   port (
      i_rst             : in std_logic
   );
end entity memory_management;

architecture rtl of memory_management is

begin



end architecture rtl;
