library ieee;
  use ieee.std_logic_1164.all;
  use IEEE.std_logic_unsigned.all;
  use IEEE.math_real.all;
  
 package select_wr_pkg is
   constant SB     : std_logic_vector(2 downto 0) := "000";
   constant SH     : std_logic_vector(2 downto 0) := "001";
   constant SW     : std_logic_vector(2 downto 0) := "010";
 end;
 
 package body select_wr_pkg is
 
 end package body;
