library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
   use ieee.numeric_std.all;
library rysy_pkg;
   use rysy_pkg.rysyPkg.all;
library ctrl_lib;
   use ctrl_lib.all;
   use ctrl_lib.ctrl_pkg.all;

entity ctrl is
   port (
   );
end entity ctrl;

architecture rtl of ctrl is


begin

   p_ctrl : process(all)
   begin

   end process p_ctrl;

end architecture rtl;
