library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
   use ieee.numeric_std.all;
library reg_file_lib;
   use reg_file_lib.all;
   use reg_file_lib.reg_file_pkg.all;

entity reg_file is
   port (
   );
end entity reg_file;

architecture rtl of reg_file is

begin

   p_reg_file : process(all)
   begin
   end process p_reg_file;

end architecture rtl;
