// SB, SH, ... are S-type instructions, storage instructions.
`define SB  3'b000
`define SH  3'b001
`define SW  3'b010
