library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
   use ieee.numeric_std.all;
library rysy_pkg;
   use rysy_pkg.rysyPkg.all;
library decode_lib;
   use decode_lib.all;
   use decode_lib.decode_pkg.all;

entity decode is
   port (
   );
end entity decode;

architecture rtl of decode is


begin

   p_decode : process(all)
   begin

   end process p_decode;

end architecture rtl;
