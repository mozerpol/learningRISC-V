library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
   use ieee.numeric_std.all;
library rysy_pkg;
   use rysy_pkg.rysyPkg.all;
library cmp_lib;
   use cmp_lib.all;
   use cmp_lib.cmp_pkg.all;

entity cmp is
   port (
   );
end entity cmp;

architecture rtl of cmp is

begin

   p_cmp : process(all)
   begin
   end process p_cmp;

end architecture rtl;
