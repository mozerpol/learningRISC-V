library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;


entity bus_interconnect is
   port (
   );
end entity bus_interconnect;

architecture rtl of bus_interconnect is

begin


end architecture rtl;
