library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
   use ieee.numeric_std.all;
library control_lib;
   use control_lib.all;
   use control_lib.control_pkg.all;

entity control is
   port (
   );
end entity control;

architecture rtl of control is

begin

   p_control : process(all)
   begin
   end process p_control;

end architecture rtl;
