library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
   use ieee.numeric_std.all;
library alu_lib;
   use alu_lib.all;
   use alu_lib.alu_pkg.all;

entity alu is
   port (
   );
end entity alu;

architecture rtl of alu is

begin

   p_alu : process(all)
   begin
   end process p_alu;

end architecture rtl;
