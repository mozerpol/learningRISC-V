library ieee;
  use ieee.std_logic_1164.all;
  use IEEE.std_logic_unsigned.all;
  use IEEE.math_real.all;
  
 package alu1_mux_pkg is
    -- constant C_NAME : std_logic_vector(N downto M) := "X";
    constant ALU1_RS   : std_logic := '0';
    constant ALU1_PC   : std_logic := '1';
 end;
 
 package body alu1_mux_pkg is
 
 end package body;
