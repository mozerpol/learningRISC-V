library ieee;
  use ieee.std_logic_1164.all;
  use IEEE.std_logic_unsigned.all;
  use IEEE.math_real.all;
  
 package byte_enabled_simple_dual_port_ram_pkg is
    -- constant C_NAME : std_logic_vector(N downto M) := "X";
    type t_array is array (integer range<>) of std_logic_vector;
 end;
 
 package body byte_enabled_simple_dual_port_ram_pkg is
 
 end package body;
