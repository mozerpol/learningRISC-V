library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;


entity byte_enabled_simple_dual_port_ram is
   port (
   );
end entity byte_enabled_simple_dual_port_ram;

architecture rtl of byte_enabled_simple_dual_port_ram is

begin


end architecture rtl;
