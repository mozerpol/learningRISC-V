`define ALU2_RS 0
`define ALU2_IMM 1