library ieee;
   use ieee.std_logic_1164.all;
   use IEEE.std_logic_unsigned.all;
   use IEEE.math_real.all;

package main_pkg is

   constant C_RAM_LENGTH      : integer := 64;
   constant C_ROM_LENGTH      : integer := 1024;
   constant C_MMIO_ADDR_GPIO  : integer := 64;

end;

package body main_pkg is

end package body;
