library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
   use ieee.numeric_std.all;
library core_lib;
   use core_lib.all;
   use core_lib.core_pkg.all;
   
   
entity core is
   port (

   );
end entity core;

architecture rtl of core is






begin





end architecture rtl;
