library ieee;
  use ieee.std_logic_1164.all;
  use IEEE.std_logic_unsigned.all;
  use IEEE.math_real.all;
  
 package alu2_mux_pkg is
    -- constant C_NAME : std_logic_vector(N downto M) := "X";
 end;
 
 package body alu2_mux_pkg is
 
 end package body;
