`define RD_IMM 	2'b00
`define RD_PCP4 	2'b01
`define RD_ALU 	2'b10
`define RD_MEM 	2'b11