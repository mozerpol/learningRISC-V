/*-
 * SPDX-License-Identifier: BSD-3-Clause
 *
 * Copyright (c) 2019 Rafal Kozik
 * All rights reserved.
 */

package selectPkg;
	typedef enum bit [2:0] {
		SB,
		SH,
		SW,
		SBU,
		SHU
	} sel_type;
endpackage : selectPkg
