library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
   use ieee.numeric_std.all;
library memory_lib;
   use memory_lib.all;
   use memory_lib.memory_pkg.all;

entity memory is
   port (
   );
end entity memory;

architecture rtl of memory is

begin

   p_memory : process(all)
   begin
   end process p_memory;

end architecture rtl;
