library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;

package rysyPkg is
   constant REG_LEN     : integer := 32;
   constant REG_NUM     : integer := 32;
   constant ADDR_LEN    : integer := 5;
   constant NOP         : integer := 13;
end;

package body rysyPkg is

end package body;
