library ieee;
  use ieee.std_logic_1164.all;
  use IEEE.std_logic_unsigned.all;
  use IEEE.math_real.all;
  
 package control_pkg is


   
 end;
 
 package body control_pkg is
 
 end package body;
