library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
library rysy_pkg;
   use rysy_pkg.rysyPkg.all;


entity reg_file_design is
   port (
   );
end entity reg_file_design;

architecture rtl of reg_file_design is

begin

end architecture rtl;
