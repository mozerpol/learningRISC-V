library ieee;
   use ieee.std_logic_1164.all;
   use ieee.numeric_std.all;
   use ieee.std_logic_unsigned.all;
library rysy_pkg;
   use rysy_pkg.rysyPkg.all;
library std;
  use std.env.all;

entity cmp_tb is
end cmp_tb;

architecture tb of cmp_tb is

   component cmp is
   port (
   );
   end component cmp;
 
begin

   inst_cmp : component cmp 
   port map (
   );

   p_tb : process
   begin
       
      wait for 25 ns;
      stop(2); 
   end process p_tb;

end architecture tb;
