`define REG_LEN 32
`define REG_NUM 32
