library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
library rysy_pkg;
   use rysy_pkg.rysyPkg.all;


entity rd_mux_design is
   port (
   );
end entity rd_mux_design;

architecture rtl of rd_mux_design is

begin

end architecture rtl;
