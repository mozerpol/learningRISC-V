`define REG_LEN 32
`define REG_NUM 32
`define ADDR_LEN 5
