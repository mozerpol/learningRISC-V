`define ALU1_RS 1'b0
`define ALU1_PC 1'b1