library ieee;
   use ieee.std_logic_1164.all;


entity alu1_mux_design is
   port (
      input rs1_d : std_logic
   );
end entity alu1_mux_design;



