library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;


entity gpio is
   port (
   );
end entity gpio;

architecture rtl of gpio is

begin


end architecture rtl;
