library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;


entity bus_interconnect_design is
   port (
   );
end entity bus_interconnect_design;

architecture rtl of bus_interconnect_design is

begin


end architecture rtl;
