library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
   use ieee.numeric_std.all;
library decoder_lib;
   use decoder_lib.all;
   use decoder_lib.decoder_pkg.all;

entity decoder is
   port (
   );
end entity decoder;

architecture rtl of decoder is

begin

   p_decoder : process(all)
   begin
   end process p_decoder;

end architecture rtl;
