library ieee;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_unsigned.all;
   use ieee.numeric_std.all;
library rysy_pkg;
   use rysy_pkg.rysyPkg.all;
library inst_mgmt_lib;
   use inst_mgmt_lib.all;
   use inst_mgmt_lib.inst_mgmt_pkg.all;

entity inst_mgmt is
   port (
   );
end entity inst_mgmt;

architecture rtl of inst_mgmt is

begin

   p_inst_mgmt : process(all)
   begin
   end process p_inst_mgmt;

end architecture rtl;
