`define REG_LEN 32
