library ieee;
   use ieee.std_logic_1164.all;
   use ieee.numeric_std.all;
   use ieee.std_logic_unsigned.all;
   
entity rysy is
   port (
      clk      : in std_logic
   );
end entity rysy;

architecture rtl of rysy is


begin

   p_rysy : process(clk)
   begin
   end process p_rysy;


end architecture rtl;
